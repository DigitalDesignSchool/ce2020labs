// y(t) = sin(2*pi*F*t), F=261.63Hz, Fs=48000Hz, 16-bit

module lut_C
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 182;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010001100101;
        2: y = 16'b0000100011001000;
        3: y = 16'b0000110100101001;
        4: y = 16'b0001000110000110;
        5: y = 16'b0001010111011110;
        6: y = 16'b0001101000101111;
        7: y = 16'b0001111001111000;
        8: y = 16'b0010001010111000;
        9: y = 16'b0010011011101101;
        10: y = 16'b0010101100010111;
        11: y = 16'b0010111100110011;
        12: y = 16'b0011001101000010;
        13: y = 16'b0011011101000001;
        14: y = 16'b0011101100101111;
        15: y = 16'b0011111100001011;
        16: y = 16'b0100001011010101;
        17: y = 16'b0100011010001010;
        18: y = 16'b0100101000101010;
        19: y = 16'b0100110110110011;
        20: y = 16'b0101000100100110;
        21: y = 16'b0101010001111111;
        22: y = 16'b0101011110111111;
        23: y = 16'b0101101011100101;
        24: y = 16'b0101110111101111;
        25: y = 16'b0110000011011101;
        26: y = 16'b0110001110101110;
        27: y = 16'b0110011001100000;
        28: y = 16'b0110100011110100;
        29: y = 16'b0110101101101000;
        30: y = 16'b0110110110111100;
        31: y = 16'b0110111111101110;
        32: y = 16'b0111000111111111;
        33: y = 16'b0111001111101101;
        34: y = 16'b0111010110111000;
        35: y = 16'b0111011101100000;
        36: y = 16'b0111100011100100;
        37: y = 16'b0111101001000011;
        38: y = 16'b0111101101111110;
        39: y = 16'b0111110010010011;
        40: y = 16'b0111110110000011;
        41: y = 16'b0111111001001100;
        42: y = 16'b0111111011110000;
        43: y = 16'b0111111101101101;
        44: y = 16'b0111111111000100;
        45: y = 16'b0111111111110100;
        46: y = 16'b0111111111111110;
        47: y = 16'b0111111111100001;
        48: y = 16'b0111111110011101;
        49: y = 16'b0111111100110011;
        50: y = 16'b0111111010100011;
        51: y = 16'b0111110111101100;
        52: y = 16'b0111110100001111;
        53: y = 16'b0111110000001101;
        54: y = 16'b0111101011100101;
        55: y = 16'b0111100110011000;
        56: y = 16'b0111100000100111;
        57: y = 16'b0111011010010001;
        58: y = 16'b0111010011010111;
        59: y = 16'b0111001011111010;
        60: y = 16'b0111000011111011;
        61: y = 16'b0110111011011001;
        62: y = 16'b0110110010010110;
        63: y = 16'b0110101000110010;
        64: y = 16'b0110011110101110;
        65: y = 16'b0110010100001011;
        66: y = 16'b0110001001001001;
        67: y = 16'b0101111101101010;
        68: y = 16'b0101110001101110;
        69: y = 16'b0101100101010110;
        70: y = 16'b0101011000100011;
        71: y = 16'b0101001011010110;
        72: y = 16'b0100111101110000;
        73: y = 16'b0100101111110010;
        74: y = 16'b0100100001011101;
        75: y = 16'b0100010010110010;
        76: y = 16'b0100000011110010;
        77: y = 16'b0011110100011111;
        78: y = 16'b0011100100111010;
        79: y = 16'b0011010101000011;
        80: y = 16'b0011000100111100;
        81: y = 16'b0010110100100111;
        82: y = 16'b0010100100000011;
        83: y = 16'b0010010011010100;
        84: y = 16'b0010000010011001;
        85: y = 16'b0001110001010100;
        86: y = 16'b0001100000000111;
        87: y = 16'b0001001110110011;
        88: y = 16'b0000111101011000;
        89: y = 16'b0000101011111001;
        90: y = 16'b0000011010010111;
        91: y = 16'b0000001000110010;
        92: y = 16'b1111110111001110;
        93: y = 16'b1111100101101001;
        94: y = 16'b1111010100000111;
        95: y = 16'b1111000010101000;
        96: y = 16'b1110110001001101;
        97: y = 16'b1110011111111001;
        98: y = 16'b1110001110101100;
        99: y = 16'b1101111101100111;
        100: y = 16'b1101101100101100;
        101: y = 16'b1101011011111101;
        102: y = 16'b1101001011011001;
        103: y = 16'b1100111011000100;
        104: y = 16'b1100101010111101;
        105: y = 16'b1100011011000110;
        106: y = 16'b1100001011100001;
        107: y = 16'b1011111100001110;
        108: y = 16'b1011101101001110;
        109: y = 16'b1011011110100011;
        110: y = 16'b1011010000001110;
        111: y = 16'b1011000010010000;
        112: y = 16'b1010110100101010;
        113: y = 16'b1010100111011101;
        114: y = 16'b1010011010101010;
        115: y = 16'b1010001110010010;
        116: y = 16'b1010000010010110;
        117: y = 16'b1001110110110111;
        118: y = 16'b1001101011110101;
        119: y = 16'b1001100001010010;
        120: y = 16'b1001010111001110;
        121: y = 16'b1001001101101010;
        122: y = 16'b1001000100100111;
        123: y = 16'b1000111100000101;
        124: y = 16'b1000110100000110;
        125: y = 16'b1000101100101001;
        126: y = 16'b1000100101101111;
        127: y = 16'b1000011111011001;
        128: y = 16'b1000011001101000;
        129: y = 16'b1000010100011011;
        130: y = 16'b1000001111110011;
        131: y = 16'b1000001011110001;
        132: y = 16'b1000001000010100;
        133: y = 16'b1000000101011101;
        134: y = 16'b1000000011001101;
        135: y = 16'b1000000001100011;
        136: y = 16'b1000000000011111;
        137: y = 16'b1000000000000010;
        138: y = 16'b1000000000001100;
        139: y = 16'b1000000000111100;
        140: y = 16'b1000000010010011;
        141: y = 16'b1000000100010000;
        142: y = 16'b1000000110110100;
        143: y = 16'b1000001001111101;
        144: y = 16'b1000001101101101;
        145: y = 16'b1000010010000010;
        146: y = 16'b1000010110111101;
        147: y = 16'b1000011100011100;
        148: y = 16'b1000100010100000;
        149: y = 16'b1000101001001000;
        150: y = 16'b1000110000010011;
        151: y = 16'b1000111000000001;
        152: y = 16'b1001000000010010;
        153: y = 16'b1001001001000100;
        154: y = 16'b1001010010011000;
        155: y = 16'b1001011100001100;
        156: y = 16'b1001100110100000;
        157: y = 16'b1001110001010010;
        158: y = 16'b1001111100100011;
        159: y = 16'b1010001000010001;
        160: y = 16'b1010010100011011;
        161: y = 16'b1010100001000001;
        162: y = 16'b1010101110000001;
        163: y = 16'b1010111011011010;
        164: y = 16'b1011001001001101;
        165: y = 16'b1011010111010110;
        166: y = 16'b1011100101110110;
        167: y = 16'b1011110100101011;
        168: y = 16'b1100000011110101;
        169: y = 16'b1100010011010001;
        170: y = 16'b1100100010111111;
        171: y = 16'b1100110010111110;
        172: y = 16'b1101000011001101;
        173: y = 16'b1101010011101001;
        174: y = 16'b1101100100010011;
        175: y = 16'b1101110101001000;
        176: y = 16'b1110000110001000;
        177: y = 16'b1110010111010001;
        178: y = 16'b1110101000100010;
        179: y = 16'b1110111001111010;
        180: y = 16'b1111001011010111;
        181: y = 16'b1111011100111000;
        182: y = 16'b1111101110011011;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=277.18Hz, Fs=48000Hz, 16-bit

module lut_Cs
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 172;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010010100110;
        2: y = 16'b0000100101001010;
        3: y = 16'b0000110111101011;
        4: y = 16'b0001001010001000;
        5: y = 16'b0001011100011110;
        6: y = 16'b0001101110101100;
        7: y = 16'b0010000000110001;
        8: y = 16'b0010010010101011;
        9: y = 16'b0010100100011001;
        10: y = 16'b0010110101111001;
        11: y = 16'b0011000111001001;
        12: y = 16'b0011011000001001;
        13: y = 16'b0011101000110110;
        14: y = 16'b0011111001010000;
        15: y = 16'b0100001001010101;
        16: y = 16'b0100011001000011;
        17: y = 16'b0100101000011010;
        18: y = 16'b0100110111011000;
        19: y = 16'b0101000101111011;
        20: y = 16'b0101010100000011;
        21: y = 16'b0101100001101110;
        22: y = 16'b0101101110111011;
        23: y = 16'b0101111011101001;
        24: y = 16'b0110000111111000;
        25: y = 16'b0110010011100101;
        26: y = 16'b0110011110110000;
        27: y = 16'b0110101001011000;
        28: y = 16'b0110110011011100;
        29: y = 16'b0110111100111100;
        30: y = 16'b0111000101110110;
        31: y = 16'b0111001110001001;
        32: y = 16'b0111010101110110;
        33: y = 16'b0111011100111011;
        34: y = 16'b0111100011010111;
        35: y = 16'b0111101001001011;
        36: y = 16'b0111101110010110;
        37: y = 16'b0111110010110110;
        38: y = 16'b0111110110101101;
        39: y = 16'b0111111001111001;
        40: y = 16'b0111111100011011;
        41: y = 16'b0111111110010010;
        42: y = 16'b0111111111011101;
        43: y = 16'b0111111111111110;
        44: y = 16'b0111111111110011;
        45: y = 16'b0111111110111101;
        46: y = 16'b0111111101011100;
        47: y = 16'b0111111011010000;
        48: y = 16'b0111111000011001;
        49: y = 16'b0111110100110111;
        50: y = 16'b0111110000101011;
        51: y = 16'b0111101011110110;
        52: y = 16'b0111100110010110;
        53: y = 16'b0111100000001110;
        54: y = 16'b0111011001011101;
        55: y = 16'b0111010010000100;
        56: y = 16'b0111001010000100;
        57: y = 16'b0111000001011101;
        58: y = 16'b0110111000010001;
        59: y = 16'b0110101110011111;
        60: y = 16'b0110100100001000;
        61: y = 16'b0110011001001111;
        62: y = 16'b0110001101110010;
        63: y = 16'b0110000001110101;
        64: y = 16'b0101110101010110;
        65: y = 16'b0101101000011000;
        66: y = 16'b0101011010111100;
        67: y = 16'b0101001101000010;
        68: y = 16'b0100111110101101;
        69: y = 16'b0100101111111100;
        70: y = 16'b0100100000110010;
        71: y = 16'b0100010001001111;
        72: y = 16'b0100000001010101;
        73: y = 16'b0011110001000110;
        74: y = 16'b0011100000100010;
        75: y = 16'b0011001111101011;
        76: y = 16'b0010111110100011;
        77: y = 16'b0010101101001011;
        78: y = 16'b0010011011100100;
        79: y = 16'b0010001001110000;
        80: y = 16'b0001110111110000;
        81: y = 16'b0001100101100110;
        82: y = 16'b0001010011010011;
        83: y = 16'b0001000000111010;
        84: y = 16'b0000101110011011;
        85: y = 16'b0000011011111000;
        86: y = 16'b0000001001010011;
        87: y = 16'b1111110110101101;
        88: y = 16'b1111100100001000;
        89: y = 16'b1111010001100101;
        90: y = 16'b1110111111000110;
        91: y = 16'b1110101100101101;
        92: y = 16'b1110011010011010;
        93: y = 16'b1110001000010000;
        94: y = 16'b1101110110010000;
        95: y = 16'b1101100100011100;
        96: y = 16'b1101010010110101;
        97: y = 16'b1101000001011101;
        98: y = 16'b1100110000010101;
        99: y = 16'b1100011111011110;
        100: y = 16'b1100001110111010;
        101: y = 16'b1011111110101011;
        102: y = 16'b1011101110110001;
        103: y = 16'b1011011111001110;
        104: y = 16'b1011010000000100;
        105: y = 16'b1011000001010011;
        106: y = 16'b1010110010111110;
        107: y = 16'b1010100101000100;
        108: y = 16'b1010010111101000;
        109: y = 16'b1010001010101010;
        110: y = 16'b1001111110001011;
        111: y = 16'b1001110010001110;
        112: y = 16'b1001100110110001;
        113: y = 16'b1001011011111000;
        114: y = 16'b1001010001100001;
        115: y = 16'b1001000111101111;
        116: y = 16'b1000111110100011;
        117: y = 16'b1000110101111100;
        118: y = 16'b1000101101111100;
        119: y = 16'b1000100110100011;
        120: y = 16'b1000011111110010;
        121: y = 16'b1000011001101010;
        122: y = 16'b1000010100001010;
        123: y = 16'b1000001111010101;
        124: y = 16'b1000001011001001;
        125: y = 16'b1000000111100111;
        126: y = 16'b1000000100110000;
        127: y = 16'b1000000010100100;
        128: y = 16'b1000000001000011;
        129: y = 16'b1000000000001101;
        130: y = 16'b1000000000000010;
        131: y = 16'b1000000000100011;
        132: y = 16'b1000000001101110;
        133: y = 16'b1000000011100101;
        134: y = 16'b1000000110000111;
        135: y = 16'b1000001001010011;
        136: y = 16'b1000001101001010;
        137: y = 16'b1000010001101010;
        138: y = 16'b1000010110110101;
        139: y = 16'b1000011100101001;
        140: y = 16'b1000100011000101;
        141: y = 16'b1000101010001010;
        142: y = 16'b1000110001110111;
        143: y = 16'b1000111010001010;
        144: y = 16'b1001000011000100;
        145: y = 16'b1001001100100100;
        146: y = 16'b1001010110101000;
        147: y = 16'b1001100001010000;
        148: y = 16'b1001101100011011;
        149: y = 16'b1001111000001000;
        150: y = 16'b1010000100010111;
        151: y = 16'b1010010001000101;
        152: y = 16'b1010011110010010;
        153: y = 16'b1010101011111101;
        154: y = 16'b1010111010000101;
        155: y = 16'b1011001000101000;
        156: y = 16'b1011010111100110;
        157: y = 16'b1011100110111101;
        158: y = 16'b1011110110101011;
        159: y = 16'b1100000110110000;
        160: y = 16'b1100010111001010;
        161: y = 16'b1100100111110111;
        162: y = 16'b1100111000110111;
        163: y = 16'b1101001010000111;
        164: y = 16'b1101011011100111;
        165: y = 16'b1101101101010101;
        166: y = 16'b1101111111001111;
        167: y = 16'b1110010001010100;
        168: y = 16'b1110100011100010;
        169: y = 16'b1110110101111000;
        170: y = 16'b1111001000010101;
        171: y = 16'b1111011010110110;
        172: y = 16'b1111101101011010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=293.66Hz, Fs=48000Hz, 16-bit

module lut_D
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 162;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010011101111;
        2: y = 16'b0000100111011100;
        3: y = 16'b0000111011000101;
        4: y = 16'b0001001110101000;
        5: y = 16'b0001100010000100;
        6: y = 16'b0001110101010111;
        7: y = 16'b0010001000011111;
        8: y = 16'b0010011011011001;
        9: y = 16'b0010101110000101;
        10: y = 16'b0011000000100000;
        11: y = 16'b0011010010101001;
        12: y = 16'b0011100100011110;
        13: y = 16'b0011110101111101;
        14: y = 16'b0100000111000101;
        15: y = 16'b0100010111110100;
        16: y = 16'b0100101000001000;
        17: y = 16'b0100111000000000;
        18: y = 16'b0101000111011011;
        19: y = 16'b0101010110010110;
        20: y = 16'b0101100100110000;
        21: y = 16'b0101110010101001;
        22: y = 16'b0101111111111111;
        23: y = 16'b0110001100110000;
        24: y = 16'b0110011000111011;
        25: y = 16'b0110100100011111;
        26: y = 16'b0110101111011100;
        27: y = 16'b0110111001101111;
        28: y = 16'b0111000011011001;
        29: y = 16'b0111001100010111;
        30: y = 16'b0111010100101010;
        31: y = 16'b0111011100010000;
        32: y = 16'b0111100011001001;
        33: y = 16'b0111101001010100;
        34: y = 16'b0111101110110000;
        35: y = 16'b0111110011011101;
        36: y = 16'b0111110111011011;
        37: y = 16'b0111111010101001;
        38: y = 16'b0111111101000111;
        39: y = 16'b0111111110110100;
        40: y = 16'b0111111111110001;
        41: y = 16'b0111111111111101;
        42: y = 16'b0111111111011001;
        43: y = 16'b0111111110000100;
        44: y = 16'b0111111011111110;
        45: y = 16'b0111111001001000;
        46: y = 16'b0111110101100010;
        47: y = 16'b0111110001001101;
        48: y = 16'b0111101100001000;
        49: y = 16'b0111100110010100;
        50: y = 16'b0111011111110010;
        51: y = 16'b0111011000100010;
        52: y = 16'b0111010000100110;
        53: y = 16'b0111000111111101;
        54: y = 16'b0110111110101001;
        55: y = 16'b0110110100101011;
        56: y = 16'b0110101010000011;
        57: y = 16'b0110011110110010;
        58: y = 16'b0110010010111010;
        59: y = 16'b0110000110011100;
        60: y = 16'b0101111001011000;
        61: y = 16'b0101101011110001;
        62: y = 16'b0101011101100111;
        63: y = 16'b0101001110111100;
        64: y = 16'b0100111111110001;
        65: y = 16'b0100110000001000;
        66: y = 16'b0100100000000001;
        67: y = 16'b0100001111100000;
        68: y = 16'b0011111110100100;
        69: y = 16'b0011101101010001;
        70: y = 16'b0011011011100110;
        71: y = 16'b0011001001100111;
        72: y = 16'b0010110111010101;
        73: y = 16'b0010100100110001;
        74: y = 16'b0010010001111110;
        75: y = 16'b0001111110111100;
        76: y = 16'b0001101011101111;
        77: y = 16'b0001011000010111;
        78: y = 16'b0001000100110111;
        79: y = 16'b0000110001010001;
        80: y = 16'b0000011101100110;
        81: y = 16'b0000001001110111;
        82: y = 16'b1111110110001001;
        83: y = 16'b1111100010011010;
        84: y = 16'b1111001110101111;
        85: y = 16'b1110111011001001;
        86: y = 16'b1110100111101001;
        87: y = 16'b1110010100010001;
        88: y = 16'b1110000001000100;
        89: y = 16'b1101101110000010;
        90: y = 16'b1101011011001111;
        91: y = 16'b1101001000101011;
        92: y = 16'b1100110110011001;
        93: y = 16'b1100100100011010;
        94: y = 16'b1100010010101111;
        95: y = 16'b1100000001011100;
        96: y = 16'b1011110000100000;
        97: y = 16'b1011011111111111;
        98: y = 16'b1011001111111000;
        99: y = 16'b1011000000001111;
        100: y = 16'b1010110001000100;
        101: y = 16'b1010100010011001;
        102: y = 16'b1010010100001111;
        103: y = 16'b1010000110101000;
        104: y = 16'b1001111001100100;
        105: y = 16'b1001101101000110;
        106: y = 16'b1001100001001110;
        107: y = 16'b1001010101111101;
        108: y = 16'b1001001011010101;
        109: y = 16'b1001000001010111;
        110: y = 16'b1000111000000011;
        111: y = 16'b1000101111011010;
        112: y = 16'b1000100111011110;
        113: y = 16'b1000100000001110;
        114: y = 16'b1000011001101100;
        115: y = 16'b1000010011111000;
        116: y = 16'b1000001110110011;
        117: y = 16'b1000001010011110;
        118: y = 16'b1000000110111000;
        119: y = 16'b1000000100000010;
        120: y = 16'b1000000001111100;
        121: y = 16'b1000000000100111;
        122: y = 16'b1000000000000011;
        123: y = 16'b1000000000001111;
        124: y = 16'b1000000001001100;
        125: y = 16'b1000000010111001;
        126: y = 16'b1000000101010111;
        127: y = 16'b1000001000100101;
        128: y = 16'b1000001100100011;
        129: y = 16'b1000010001010000;
        130: y = 16'b1000010110101100;
        131: y = 16'b1000011100110111;
        132: y = 16'b1000100011110000;
        133: y = 16'b1000101011010110;
        134: y = 16'b1000110011101001;
        135: y = 16'b1000111100100111;
        136: y = 16'b1001000110010001;
        137: y = 16'b1001010000100100;
        138: y = 16'b1001011011100001;
        139: y = 16'b1001100111000101;
        140: y = 16'b1001110011010000;
        141: y = 16'b1010000000000001;
        142: y = 16'b1010001101010111;
        143: y = 16'b1010011011010000;
        144: y = 16'b1010101001101010;
        145: y = 16'b1010111000100101;
        146: y = 16'b1011001000000000;
        147: y = 16'b1011010111111000;
        148: y = 16'b1011101000001100;
        149: y = 16'b1011111000111011;
        150: y = 16'b1100001010000011;
        151: y = 16'b1100011011100010;
        152: y = 16'b1100101101010111;
        153: y = 16'b1100111111100000;
        154: y = 16'b1101010001111011;
        155: y = 16'b1101100100100111;
        156: y = 16'b1101110111100001;
        157: y = 16'b1110001010101001;
        158: y = 16'b1110011101111100;
        159: y = 16'b1110110001011000;
        160: y = 16'b1111000100111011;
        161: y = 16'b1111011000100100;
        162: y = 16'b1111101100010001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=311.13Hz, Fs=48000Hz, 16-bit

module lut_Ds
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 153;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010100111001;
        2: y = 16'b0000101001101111;
        3: y = 16'b0000111110100001;
        4: y = 16'b0001010011001100;
        5: y = 16'b0001100111101110;
        6: y = 16'b0001111100000101;
        7: y = 16'b0010010000010000;
        8: y = 16'b0010100100001010;
        9: y = 16'b0010110111110011;
        10: y = 16'b0011001011001001;
        11: y = 16'b0011011110001001;
        12: y = 16'b0011110000110001;
        13: y = 16'b0100000011000000;
        14: y = 16'b0100010100110011;
        15: y = 16'b0100100110001001;
        16: y = 16'b0100110110111111;
        17: y = 16'b0101000111010100;
        18: y = 16'b0101010111000110;
        19: y = 16'b0101100110010100;
        20: y = 16'b0101110100111100;
        21: y = 16'b0110000010111100;
        22: y = 16'b0110010000010010;
        23: y = 16'b0110011100111110;
        24: y = 16'b0110101000111110;
        25: y = 16'b0110110100010001;
        26: y = 16'b0110111110110101;
        27: y = 16'b0111001000101010;
        28: y = 16'b0111010001101110;
        29: y = 16'b0111011010000000;
        30: y = 16'b0111100001100000;
        31: y = 16'b0111101000001101;
        32: y = 16'b0111101110000101;
        33: y = 16'b0111110011001001;
        34: y = 16'b0111110111011000;
        35: y = 16'b0111111010110001;
        36: y = 16'b0111111101010101;
        37: y = 16'b0111111111000010;
        38: y = 16'b0111111111111000;
        39: y = 16'b0111111111111000;
        40: y = 16'b0111111111000010;
        41: y = 16'b0111111101010101;
        42: y = 16'b0111111010110001;
        43: y = 16'b0111110111011000;
        44: y = 16'b0111110011001001;
        45: y = 16'b0111101110000101;
        46: y = 16'b0111101000001101;
        47: y = 16'b0111100001100000;
        48: y = 16'b0111011010000000;
        49: y = 16'b0111010001101110;
        50: y = 16'b0111001000101010;
        51: y = 16'b0110111110110101;
        52: y = 16'b0110110100010001;
        53: y = 16'b0110101000111110;
        54: y = 16'b0110011100111110;
        55: y = 16'b0110010000010010;
        56: y = 16'b0110000010111100;
        57: y = 16'b0101110100111100;
        58: y = 16'b0101100110010100;
        59: y = 16'b0101010111000110;
        60: y = 16'b0101000111010100;
        61: y = 16'b0100110110111111;
        62: y = 16'b0100100110001001;
        63: y = 16'b0100010100110011;
        64: y = 16'b0100000011000000;
        65: y = 16'b0011110000110001;
        66: y = 16'b0011011110001001;
        67: y = 16'b0011001011001001;
        68: y = 16'b0010110111110011;
        69: y = 16'b0010100100001010;
        70: y = 16'b0010010000010000;
        71: y = 16'b0001111100000101;
        72: y = 16'b0001100111101110;
        73: y = 16'b0001010011001100;
        74: y = 16'b0000111110100001;
        75: y = 16'b0000101001101111;
        76: y = 16'b0000010100111001;
        77: y = 16'b0000000000000000;
        78: y = 16'b1111101011000111;
        79: y = 16'b1111010110010001;
        80: y = 16'b1111000001011111;
        81: y = 16'b1110101100110100;
        82: y = 16'b1110011000010010;
        83: y = 16'b1110000011111011;
        84: y = 16'b1101101111110000;
        85: y = 16'b1101011011110110;
        86: y = 16'b1101001000001101;
        87: y = 16'b1100110100110111;
        88: y = 16'b1100100001110111;
        89: y = 16'b1100001111001111;
        90: y = 16'b1011111101000000;
        91: y = 16'b1011101011001101;
        92: y = 16'b1011011001110111;
        93: y = 16'b1011001001000001;
        94: y = 16'b1010111000101100;
        95: y = 16'b1010101000111010;
        96: y = 16'b1010011001101100;
        97: y = 16'b1010001011000100;
        98: y = 16'b1001111101000100;
        99: y = 16'b1001101111101110;
        100: y = 16'b1001100011000010;
        101: y = 16'b1001010111000010;
        102: y = 16'b1001001011101111;
        103: y = 16'b1001000001001011;
        104: y = 16'b1000110111010110;
        105: y = 16'b1000101110010010;
        106: y = 16'b1000100110000000;
        107: y = 16'b1000011110100000;
        108: y = 16'b1000010111110011;
        109: y = 16'b1000010001111011;
        110: y = 16'b1000001100110111;
        111: y = 16'b1000001000101000;
        112: y = 16'b1000000101001111;
        113: y = 16'b1000000010101011;
        114: y = 16'b1000000000111110;
        115: y = 16'b1000000000001000;
        116: y = 16'b1000000000001000;
        117: y = 16'b1000000000111110;
        118: y = 16'b1000000010101011;
        119: y = 16'b1000000101001111;
        120: y = 16'b1000001000101000;
        121: y = 16'b1000001100110111;
        122: y = 16'b1000010001111011;
        123: y = 16'b1000010111110011;
        124: y = 16'b1000011110100000;
        125: y = 16'b1000100110000000;
        126: y = 16'b1000101110010010;
        127: y = 16'b1000110111010110;
        128: y = 16'b1001000001001011;
        129: y = 16'b1001001011101111;
        130: y = 16'b1001010111000010;
        131: y = 16'b1001100011000010;
        132: y = 16'b1001101111101110;
        133: y = 16'b1001111101000100;
        134: y = 16'b1010001011000100;
        135: y = 16'b1010011001101100;
        136: y = 16'b1010101000111010;
        137: y = 16'b1010111000101100;
        138: y = 16'b1011001001000001;
        139: y = 16'b1011011001110111;
        140: y = 16'b1011101011001101;
        141: y = 16'b1011111101000000;
        142: y = 16'b1100001111001111;
        143: y = 16'b1100100001110111;
        144: y = 16'b1100110100110111;
        145: y = 16'b1101001000001101;
        146: y = 16'b1101011011110110;
        147: y = 16'b1101101111110000;
        148: y = 16'b1110000011111011;
        149: y = 16'b1110011000010010;
        150: y = 16'b1110101100110100;
        151: y = 16'b1111000001011111;
        152: y = 16'b1111010110010001;
        153: y = 16'b1111101011000111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=329.63Hz, Fs=48000Hz, 16-bit

module lut_E
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 144;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010110001011;
        2: y = 16'b0000101100010100;
        3: y = 16'b0001000010011000;
        4: y = 16'b0001011000010011;
        5: y = 16'b0001101110000100;
        6: y = 16'b0010000011101000;
        7: y = 16'b0010011000111011;
        8: y = 16'b0010101101111101;
        9: y = 16'b0011000010101001;
        10: y = 16'b0011010110111111;
        11: y = 16'b0011101010111010;
        12: y = 16'b0011111110011001;
        13: y = 16'b0100010001011001;
        14: y = 16'b0100100011111001;
        15: y = 16'b0100110101110110;
        16: y = 16'b0101000111001101;
        17: y = 16'b0101010111111101;
        18: y = 16'b0101101000000100;
        19: y = 16'b0101110111011111;
        20: y = 16'b0110000110001110;
        21: y = 16'b0110010100001101;
        22: y = 16'b0110100001011100;
        23: y = 16'b0110101101111001;
        24: y = 16'b0110111001100010;
        25: y = 16'b0111000100010110;
        26: y = 16'b0111001110010100;
        27: y = 16'b0111010111011010;
        28: y = 16'b0111011111100111;
        29: y = 16'b0111100110111011;
        30: y = 16'b0111101101010101;
        31: y = 16'b0111110010110011;
        32: y = 16'b0111110111010101;
        33: y = 16'b0111111010111011;
        34: y = 16'b0111111101100011;
        35: y = 16'b0111111111001111;
        36: y = 16'b0111111111111101;
        37: y = 16'b0111111111101110;
        38: y = 16'b0111111110100001;
        39: y = 16'b0111111100010111;
        40: y = 16'b0111111001001111;
        41: y = 16'b0111110101001011;
        42: y = 16'b0111110000001011;
        43: y = 16'b0111101010001111;
        44: y = 16'b0111100011011001;
        45: y = 16'b0111011011101000;
        46: y = 16'b0111010010111110;
        47: y = 16'b0111001001011100;
        48: y = 16'b0110111111000011;
        49: y = 16'b0110110011110100;
        50: y = 16'b0110100111110001;
        51: y = 16'b0110011010111011;
        52: y = 16'b0110001101010011;
        53: y = 16'b0101111110111100;
        54: y = 16'b0101101111110111;
        55: y = 16'b0101100000000110;
        56: y = 16'b0101001111101010;
        57: y = 16'b0100111110100110;
        58: y = 16'b0100101100111100;
        59: y = 16'b0100011010101110;
        60: y = 16'b0100000111111101;
        61: y = 16'b0011110100101101;
        62: y = 16'b0011100001000000;
        63: y = 16'b0011001100110111;
        64: y = 16'b0010111000010110;
        65: y = 16'b0010100011011111;
        66: y = 16'b0010001110010100;
        67: y = 16'b0001111000111000;
        68: y = 16'b0001100011001101;
        69: y = 16'b0001001101010111;
        70: y = 16'b0000110111010111;
        71: y = 16'b0000100001010000;
        72: y = 16'b0000001011000110;
        73: y = 16'b1111110100111010;
        74: y = 16'b1111011110110000;
        75: y = 16'b1111001000101001;
        76: y = 16'b1110110010101001;
        77: y = 16'b1110011100110011;
        78: y = 16'b1110000111001000;
        79: y = 16'b1101110001101100;
        80: y = 16'b1101011100100001;
        81: y = 16'b1101000111101010;
        82: y = 16'b1100110011001001;
        83: y = 16'b1100011111000000;
        84: y = 16'b1100001011010011;
        85: y = 16'b1011111000000011;
        86: y = 16'b1011100101010010;
        87: y = 16'b1011010011000100;
        88: y = 16'b1011000001011010;
        89: y = 16'b1010110000010110;
        90: y = 16'b1010011111111010;
        91: y = 16'b1010010000001001;
        92: y = 16'b1010000001000100;
        93: y = 16'b1001110010101101;
        94: y = 16'b1001100101000101;
        95: y = 16'b1001011000001111;
        96: y = 16'b1001001100001100;
        97: y = 16'b1001000000111101;
        98: y = 16'b1000110110100100;
        99: y = 16'b1000101101000010;
        100: y = 16'b1000100100011000;
        101: y = 16'b1000011100100111;
        102: y = 16'b1000010101110001;
        103: y = 16'b1000001111110101;
        104: y = 16'b1000001010110101;
        105: y = 16'b1000000110110001;
        106: y = 16'b1000000011101001;
        107: y = 16'b1000000001011111;
        108: y = 16'b1000000000010010;
        109: y = 16'b1000000000000011;
        110: y = 16'b1000000000110001;
        111: y = 16'b1000000010011101;
        112: y = 16'b1000000101000101;
        113: y = 16'b1000001000101011;
        114: y = 16'b1000001101001101;
        115: y = 16'b1000010010101011;
        116: y = 16'b1000011001000101;
        117: y = 16'b1000100000011001;
        118: y = 16'b1000101000100110;
        119: y = 16'b1000110001101100;
        120: y = 16'b1000111011101010;
        121: y = 16'b1001000110011110;
        122: y = 16'b1001010010000111;
        123: y = 16'b1001011110100100;
        124: y = 16'b1001101011110011;
        125: y = 16'b1001111001110010;
        126: y = 16'b1010001000100001;
        127: y = 16'b1010010111111100;
        128: y = 16'b1010101000000011;
        129: y = 16'b1010111000110011;
        130: y = 16'b1011001010001010;
        131: y = 16'b1011011100000111;
        132: y = 16'b1011101110100111;
        133: y = 16'b1100000001100111;
        134: y = 16'b1100010101000110;
        135: y = 16'b1100101001000001;
        136: y = 16'b1100111101010111;
        137: y = 16'b1101010010000011;
        138: y = 16'b1101100111000101;
        139: y = 16'b1101111100011000;
        140: y = 16'b1110010001111100;
        141: y = 16'b1110100111101101;
        142: y = 16'b1110111101101000;
        143: y = 16'b1111010011101100;
        144: y = 16'b1111101001110101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=349.23Hz, Fs=48000Hz, 16-bit

module lut_F
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 136;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010111011110;
        2: y = 16'b0000101110111001;
        3: y = 16'b0001000110001110;
        4: y = 16'b0001011101011001;
        5: y = 16'b0001110100011000;
        6: y = 16'b0010001011000111;
        7: y = 16'b0010100001100100;
        8: y = 16'b0010110111101010;
        9: y = 16'b0011001101011000;
        10: y = 16'b0011100010101011;
        11: y = 16'b0011110111011110;
        12: y = 16'b0100001011110001;
        13: y = 16'b0100011111011111;
        14: y = 16'b0100110010100111;
        15: y = 16'b0101000101000101;
        16: y = 16'b0101010110111000;
        17: y = 16'b0101100111111101;
        18: y = 16'b0101111000010001;
        19: y = 16'b0110000111110010;
        20: y = 16'b0110010110011111;
        21: y = 16'b0110100100010101;
        22: y = 16'b0110110001010010;
        23: y = 16'b0110111101010101;
        24: y = 16'b0111001000011101;
        25: y = 16'b0111010010100110;
        26: y = 16'b0111011011110001;
        27: y = 16'b0111100011111100;
        28: y = 16'b0111101011000110;
        29: y = 16'b0111110001001110;
        30: y = 16'b0111110110010011;
        31: y = 16'b0111111010010100;
        32: y = 16'b0111111101010001;
        33: y = 16'b0111111111001001;
        34: y = 16'b0111111111111101;
        35: y = 16'b0111111111101100;
        36: y = 16'b0111111110010110;
        37: y = 16'b0111111011111011;
        38: y = 16'b0111111000011100;
        39: y = 16'b0111110011111001;
        40: y = 16'b0111101110010010;
        41: y = 16'b0111100111101001;
        42: y = 16'b0111011111111111;
        43: y = 16'b0111010111010100;
        44: y = 16'b0111001101101001;
        45: y = 16'b0111000011000001;
        46: y = 16'b0110110111011011;
        47: y = 16'b0110101010111011;
        48: y = 16'b0110011101100001;
        49: y = 16'b0110001111001111;
        50: y = 16'b0110000000001000;
        51: y = 16'b0101110000001101;
        52: y = 16'b0101011111100000;
        53: y = 16'b0101001110000100;
        54: y = 16'b0100111011111011;
        55: y = 16'b0100101001001000;
        56: y = 16'b0100010101101101;
        57: y = 16'b0100000001101100;
        58: y = 16'b0011101101001000;
        59: y = 16'b0011011000000101;
        60: y = 16'b0011000010100101;
        61: y = 16'b0010101100101010;
        62: y = 16'b0010010110011000;
        63: y = 16'b0001111111110010;
        64: y = 16'b0001101000111011;
        65: y = 16'b0001010001110101;
        66: y = 16'b0000111010100101;
        67: y = 16'b0000100011001100;
        68: y = 16'b0000001011101111;
        69: y = 16'b1111110100010001;
        70: y = 16'b1111011100110100;
        71: y = 16'b1111000101011011;
        72: y = 16'b1110101110001011;
        73: y = 16'b1110010111000101;
        74: y = 16'b1110000000001110;
        75: y = 16'b1101101001101000;
        76: y = 16'b1101010011010110;
        77: y = 16'b1100111101011011;
        78: y = 16'b1100100111111011;
        79: y = 16'b1100010010111000;
        80: y = 16'b1011111110010100;
        81: y = 16'b1011101010010011;
        82: y = 16'b1011010110111000;
        83: y = 16'b1011000100000101;
        84: y = 16'b1010110001111100;
        85: y = 16'b1010100000100000;
        86: y = 16'b1010001111110011;
        87: y = 16'b1001111111111000;
        88: y = 16'b1001110000110001;
        89: y = 16'b1001100010011111;
        90: y = 16'b1001010101000101;
        91: y = 16'b1001001000100101;
        92: y = 16'b1000111100111111;
        93: y = 16'b1000110010010111;
        94: y = 16'b1000101000101100;
        95: y = 16'b1000100000000001;
        96: y = 16'b1000011000010111;
        97: y = 16'b1000010001101110;
        98: y = 16'b1000001100000111;
        99: y = 16'b1000000111100100;
        100: y = 16'b1000000100000101;
        101: y = 16'b1000000001101010;
        102: y = 16'b1000000000010100;
        103: y = 16'b1000000000000011;
        104: y = 16'b1000000000110111;
        105: y = 16'b1000000010101111;
        106: y = 16'b1000000101101100;
        107: y = 16'b1000001001101101;
        108: y = 16'b1000001110110010;
        109: y = 16'b1000010100111010;
        110: y = 16'b1000011100000100;
        111: y = 16'b1000100100001111;
        112: y = 16'b1000101101011010;
        113: y = 16'b1000110111100011;
        114: y = 16'b1001000010101011;
        115: y = 16'b1001001110101110;
        116: y = 16'b1001011011101011;
        117: y = 16'b1001101001100001;
        118: y = 16'b1001111000001110;
        119: y = 16'b1010000111101111;
        120: y = 16'b1010011000000011;
        121: y = 16'b1010101001001000;
        122: y = 16'b1010111010111011;
        123: y = 16'b1011001101011001;
        124: y = 16'b1011100000100001;
        125: y = 16'b1011110100001111;
        126: y = 16'b1100001000100010;
        127: y = 16'b1100011101010101;
        128: y = 16'b1100110010101000;
        129: y = 16'b1101001000010110;
        130: y = 16'b1101011110011100;
        131: y = 16'b1101110100111001;
        132: y = 16'b1110001011101000;
        133: y = 16'b1110100010100111;
        134: y = 16'b1110111001110010;
        135: y = 16'b1111010001000111;
        136: y = 16'b1111101000100010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=369.99Hz, Fs=48000Hz, 16-bit

module lut_Fs
(
    input      [7:0] x,
    output     [7:0] x_max,
    output reg [15:0] y
);

    assign x_max = 128;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011000111011;
        2: y = 16'b0000110001110011;
        3: y = 16'b0001001010100011;
        4: y = 16'b0001100011001000;
        5: y = 16'b0001111011011101;
        6: y = 16'b0010010011100000;
        7: y = 16'b0010101011001101;
        8: y = 16'b0011000010011111;
        9: y = 16'b0011011001010100;
        10: y = 16'b0011101111101000;
        11: y = 16'b0100000101011000;
        12: y = 16'b0100011010100000;
        13: y = 16'b0100101110111101;
        14: y = 16'b0101000010101100;
        15: y = 16'b0101010101101010;
        16: y = 16'b0101100111110100;
        17: y = 16'b0101111001001000;
        18: y = 16'b0110001001100010;
        19: y = 16'b0110011001000001;
        20: y = 16'b0110100111100001;
        21: y = 16'b0110110101000010;
        22: y = 16'b0111000001100000;
        23: y = 16'b0111001100111001;
        24: y = 16'b0111010111001101;
        25: y = 16'b0111100000011001;
        26: y = 16'b0111101000011100;
        27: y = 16'b0111101111010110;
        28: y = 16'b0111110101000011;
        29: y = 16'b0111111001100101;
        30: y = 16'b0111111100111010;
        31: y = 16'b0111111111000010;
        32: y = 16'b0111111111111101;
        33: y = 16'b0111111111101001;
        34: y = 16'b0111111110001000;
        35: y = 16'b0111111011011010;
        36: y = 16'b0111110111011110;
        37: y = 16'b0111110010010110;
        38: y = 16'b0111101100000010;
        39: y = 16'b0111100100100100;
        40: y = 16'b0111011011111100;
        41: y = 16'b0111010010001100;
        42: y = 16'b0111000111010101;
        43: y = 16'b0110111011011001;
        44: y = 16'b0110101110011010;
        45: y = 16'b0110100000011001;
        46: y = 16'b0110010001011001;
        47: y = 16'b0110000001011100;
        48: y = 16'b0101110000100101;
        49: y = 16'b0101011110110110;
        50: y = 16'b0101001100010001;
        51: y = 16'b0100111000111010;
        52: y = 16'b0100100100110100;
        53: y = 16'b0100010000000001;
        54: y = 16'b0011111010100101;
        55: y = 16'b0011100100100011;
        56: y = 16'b0011001101111110;
        57: y = 16'b0010110110111001;
        58: y = 16'b0010011111011001;
        59: y = 16'b0010000111100001;
        60: y = 16'b0001101111010101;
        61: y = 16'b0001010110110111;
        62: y = 16'b0000111110001100;
        63: y = 16'b0000100101011000;
        64: y = 16'b0000001100011110;
        65: y = 16'b1111110011100010;
        66: y = 16'b1111011010101000;
        67: y = 16'b1111000001110100;
        68: y = 16'b1110101001001001;
        69: y = 16'b1110010000101011;
        70: y = 16'b1101111000011111;
        71: y = 16'b1101100000100111;
        72: y = 16'b1101001001000111;
        73: y = 16'b1100110010000010;
        74: y = 16'b1100011011011101;
        75: y = 16'b1100000101011011;
        76: y = 16'b1011101111111111;
        77: y = 16'b1011011011001100;
        78: y = 16'b1011000111000110;
        79: y = 16'b1010110011101111;
        80: y = 16'b1010100001001010;
        81: y = 16'b1010001111011011;
        82: y = 16'b1001111110100100;
        83: y = 16'b1001101110100111;
        84: y = 16'b1001011111100111;
        85: y = 16'b1001010001100110;
        86: y = 16'b1001000100100111;
        87: y = 16'b1000111000101011;
        88: y = 16'b1000101101110100;
        89: y = 16'b1000100100000100;
        90: y = 16'b1000011011011100;
        91: y = 16'b1000010011111110;
        92: y = 16'b1000001101101010;
        93: y = 16'b1000001000100010;
        94: y = 16'b1000000100100110;
        95: y = 16'b1000000001111000;
        96: y = 16'b1000000000010111;
        97: y = 16'b1000000000000011;
        98: y = 16'b1000000000111110;
        99: y = 16'b1000000011000110;
        100: y = 16'b1000000110011011;
        101: y = 16'b1000001010111101;
        102: y = 16'b1000010000101010;
        103: y = 16'b1000010111100100;
        104: y = 16'b1000011111100111;
        105: y = 16'b1000101000110011;
        106: y = 16'b1000110011000111;
        107: y = 16'b1000111110100000;
        108: y = 16'b1001001010111110;
        109: y = 16'b1001011000011111;
        110: y = 16'b1001100110111111;
        111: y = 16'b1001110110011110;
        112: y = 16'b1010000110111000;
        113: y = 16'b1010011000001100;
        114: y = 16'b1010101010010110;
        115: y = 16'b1010111101010100;
        116: y = 16'b1011010001000011;
        117: y = 16'b1011100101100000;
        118: y = 16'b1011111010101000;
        119: y = 16'b1100010000011000;
        120: y = 16'b1100100110101100;
        121: y = 16'b1100111101100001;
        122: y = 16'b1101010100110011;
        123: y = 16'b1101101100100000;
        124: y = 16'b1110000100100011;
        125: y = 16'b1110011100111000;
        126: y = 16'b1110110101011101;
        127: y = 16'b1111001110001101;
        128: y = 16'b1111100111000101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=392.0Hz, Fs=48000Hz, 16-bit

module lut_G
(
    input      [6:0] x,
    output     [6:0] x_max,
    output reg [15:0] y
);

    assign x_max = 121;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011010010111;
        2: y = 16'b0000110100101001;
        3: y = 16'b0001001110110011;
        4: y = 16'b0001101000101111;
        5: y = 16'b0010000010011001;
        6: y = 16'b0010011011101101;
        7: y = 16'b0010110100100111;
        8: y = 16'b0011001101000010;
        9: y = 16'b0011100100111010;
        10: y = 16'b0011111100001011;
        11: y = 16'b0100010010110010;
        12: y = 16'b0100101000101010;
        13: y = 16'b0100111101110000;
        14: y = 16'b0101010001111111;
        15: y = 16'b0101100101010110;
        16: y = 16'b0101110111101111;
        17: y = 16'b0110001001001001;
        18: y = 16'b0110011001100000;
        19: y = 16'b0110101000110010;
        20: y = 16'b0110110110111100;
        21: y = 16'b0111000011111011;
        22: y = 16'b0111001111101101;
        23: y = 16'b0111011010010001;
        24: y = 16'b0111100011100100;
        25: y = 16'b0111101011100101;
        26: y = 16'b0111110010010011;
        27: y = 16'b0111110111101100;
        28: y = 16'b0111111011110000;
        29: y = 16'b0111111110011101;
        30: y = 16'b0111111111110100;
        31: y = 16'b0111111111110100;
        32: y = 16'b0111111110011101;
        33: y = 16'b0111111011110000;
        34: y = 16'b0111110111101100;
        35: y = 16'b0111110010010011;
        36: y = 16'b0111101011100101;
        37: y = 16'b0111100011100100;
        38: y = 16'b0111011010010001;
        39: y = 16'b0111001111101101;
        40: y = 16'b0111000011111011;
        41: y = 16'b0110110110111100;
        42: y = 16'b0110101000110010;
        43: y = 16'b0110011001100000;
        44: y = 16'b0110001001001001;
        45: y = 16'b0101110111101111;
        46: y = 16'b0101100101010110;
        47: y = 16'b0101010001111111;
        48: y = 16'b0100111101110000;
        49: y = 16'b0100101000101010;
        50: y = 16'b0100010010110010;
        51: y = 16'b0011111100001011;
        52: y = 16'b0011100100111010;
        53: y = 16'b0011001101000010;
        54: y = 16'b0010110100100111;
        55: y = 16'b0010011011101101;
        56: y = 16'b0010000010011001;
        57: y = 16'b0001101000101111;
        58: y = 16'b0001001110110011;
        59: y = 16'b0000110100101001;
        60: y = 16'b0000011010010111;
        61: y = 16'b0000000000000000;
        62: y = 16'b1111100101101001;
        63: y = 16'b1111001011010111;
        64: y = 16'b1110110001001101;
        65: y = 16'b1110010111010001;
        66: y = 16'b1101111101100111;
        67: y = 16'b1101100100010011;
        68: y = 16'b1101001011011001;
        69: y = 16'b1100110010111110;
        70: y = 16'b1100011011000110;
        71: y = 16'b1100000011110101;
        72: y = 16'b1011101101001110;
        73: y = 16'b1011010111010110;
        74: y = 16'b1011000010010000;
        75: y = 16'b1010101110000001;
        76: y = 16'b1010011010101010;
        77: y = 16'b1010001000010001;
        78: y = 16'b1001110110110111;
        79: y = 16'b1001100110100000;
        80: y = 16'b1001010111001110;
        81: y = 16'b1001001001000100;
        82: y = 16'b1000111100000101;
        83: y = 16'b1000110000010011;
        84: y = 16'b1000100101101111;
        85: y = 16'b1000011100011100;
        86: y = 16'b1000010100011011;
        87: y = 16'b1000001101101101;
        88: y = 16'b1000001000010100;
        89: y = 16'b1000000100010000;
        90: y = 16'b1000000001100011;
        91: y = 16'b1000000000001100;
        92: y = 16'b1000000000001100;
        93: y = 16'b1000000001100011;
        94: y = 16'b1000000100010000;
        95: y = 16'b1000001000010100;
        96: y = 16'b1000001101101101;
        97: y = 16'b1000010100011011;
        98: y = 16'b1000011100011100;
        99: y = 16'b1000100101101111;
        100: y = 16'b1000110000010011;
        101: y = 16'b1000111100000101;
        102: y = 16'b1001001001000100;
        103: y = 16'b1001010111001110;
        104: y = 16'b1001100110100000;
        105: y = 16'b1001110110110111;
        106: y = 16'b1010001000010001;
        107: y = 16'b1010011010101010;
        108: y = 16'b1010101110000001;
        109: y = 16'b1011000010010000;
        110: y = 16'b1011010111010110;
        111: y = 16'b1011101101001110;
        112: y = 16'b1100000011110101;
        113: y = 16'b1100011011000110;
        114: y = 16'b1100110010111110;
        115: y = 16'b1101001011011001;
        116: y = 16'b1101100100010011;
        117: y = 16'b1101111101100111;
        118: y = 16'b1110010111010001;
        119: y = 16'b1110110001001101;
        120: y = 16'b1111001011010111;
        121: y = 16'b1111100101101001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=415.3Hz, Fs=48000Hz, 16-bit

module lut_Gs
(
    input      [6:0] x,
    output     [6:0] x_max,
    output reg [15:0] y
);

    assign x_max = 114;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011011111101;
        2: y = 16'b0000110111110101;
        3: y = 16'b0001010011100011;
        4: y = 16'b0001101111000000;
        5: y = 16'b0010001010001000;
        6: y = 16'b0010100100110110;
        7: y = 16'b0010111111000101;
        8: y = 16'b0011011000101110;
        9: y = 16'b0011110001101111;
        10: y = 16'b0100001010000001;
        11: y = 16'b0100100001100001;
        12: y = 16'b0100111000001001;
        13: y = 16'b0101001101110101;
        14: y = 16'b0101100010100010;
        15: y = 16'b0101110110001011;
        16: y = 16'b0110001000101101;
        17: y = 16'b0110011010000100;
        18: y = 16'b0110101010001100;
        19: y = 16'b0110111001000011;
        20: y = 16'b0111000110100101;
        21: y = 16'b0111010010110001;
        22: y = 16'b0111011101100100;
        23: y = 16'b0111100110111011;
        24: y = 16'b0111101110110110;
        25: y = 16'b0111110101010010;
        26: y = 16'b0111111010001110;
        27: y = 16'b0111111101101001;
        28: y = 16'b0111111111100011;
        29: y = 16'b0111111111111100;
        30: y = 16'b0111111110110011;
        31: y = 16'b0111111100001000;
        32: y = 16'b0111110111111100;
        33: y = 16'b0111110010010000;
        34: y = 16'b0111101011000100;
        35: y = 16'b0111100010011011;
        36: y = 16'b0111011000010110;
        37: y = 16'b0111001100110110;
        38: y = 16'b0110111111111111;
        39: y = 16'b0110110001110010;
        40: y = 16'b0110100010010010;
        41: y = 16'b0110010001100010;
        42: y = 16'b0101111111100101;
        43: y = 16'b0101101100011111;
        44: y = 16'b0101011000010100;
        45: y = 16'b0101000011000111;
        46: y = 16'b0100101100111100;
        47: y = 16'b0100010101111000;
        48: y = 16'b0011111101111110;
        49: y = 16'b0011100101010100;
        50: y = 16'b0011001011111110;
        51: y = 16'b0010110010000010;
        52: y = 16'b0010010111100011;
        53: y = 16'b0001111100100111;
        54: y = 16'b0001100001010100;
        55: y = 16'b0001000101101110;
        56: y = 16'b0000101001111010;
        57: y = 16'b0000001101111111;
        58: y = 16'b1111110010000001;
        59: y = 16'b1111010110000110;
        60: y = 16'b1110111010010010;
        61: y = 16'b1110011110101100;
        62: y = 16'b1110000011011001;
        63: y = 16'b1101101000011101;
        64: y = 16'b1101001101111110;
        65: y = 16'b1100110100000010;
        66: y = 16'b1100011010101100;
        67: y = 16'b1100000010000010;
        68: y = 16'b1011101010001000;
        69: y = 16'b1011010011000100;
        70: y = 16'b1010111100111001;
        71: y = 16'b1010100111101100;
        72: y = 16'b1010010011100001;
        73: y = 16'b1010000000011011;
        74: y = 16'b1001101110011110;
        75: y = 16'b1001011101101110;
        76: y = 16'b1001001110001110;
        77: y = 16'b1001000000000001;
        78: y = 16'b1000110011001010;
        79: y = 16'b1000100111101010;
        80: y = 16'b1000011101100101;
        81: y = 16'b1000010100111100;
        82: y = 16'b1000001101110000;
        83: y = 16'b1000001000000100;
        84: y = 16'b1000000011111000;
        85: y = 16'b1000000001001101;
        86: y = 16'b1000000000000100;
        87: y = 16'b1000000000011101;
        88: y = 16'b1000000010010111;
        89: y = 16'b1000000101110010;
        90: y = 16'b1000001010101110;
        91: y = 16'b1000010001001010;
        92: y = 16'b1000011001000101;
        93: y = 16'b1000100010011100;
        94: y = 16'b1000101101001111;
        95: y = 16'b1000111001011011;
        96: y = 16'b1001000110111101;
        97: y = 16'b1001010101110100;
        98: y = 16'b1001100101111100;
        99: y = 16'b1001110111010011;
        100: y = 16'b1010001001110101;
        101: y = 16'b1010011101011110;
        102: y = 16'b1010110010001011;
        103: y = 16'b1011000111110111;
        104: y = 16'b1011011110011111;
        105: y = 16'b1011110101111111;
        106: y = 16'b1100001110010001;
        107: y = 16'b1100100111010010;
        108: y = 16'b1101000000111011;
        109: y = 16'b1101011011001010;
        110: y = 16'b1101110101111000;
        111: y = 16'b1110010001000000;
        112: y = 16'b1110101100011101;
        113: y = 16'b1111001000001011;
        114: y = 16'b1111100100000011;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=440.0Hz, Fs=48000Hz, 16-bit

module lut_A
(
    input      [6:0] x,
    output     [6:0] x_max,
    output reg [15:0] y
);

    assign x_max = 108;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011101100000;
        2: y = 16'b0000111010111001;
        3: y = 16'b0001011000000110;
        4: y = 16'b0001110101000001;
        5: y = 16'b0010010001100010;
        6: y = 16'b0010101101100100;
        7: y = 16'b0011001001000010;
        8: y = 16'b0011100011110101;
        9: y = 16'b0011111101110111;
        10: y = 16'b0100010111000011;
        11: y = 16'b0100101111010100;
        12: y = 16'b0101000110100101;
        13: y = 16'b0101011100110000;
        14: y = 16'b0101110001110001;
        15: y = 16'b0110000101100100;
        16: y = 16'b0110011000000011;
        17: y = 16'b0110101001001100;
        18: y = 16'b0110111000111010;
        19: y = 16'b0111000111001011;
        20: y = 16'b0111010011111011;
        21: y = 16'b0111011111000111;
        22: y = 16'b0111101000101110;
        23: y = 16'b0111110000101101;
        24: y = 16'b0111110111000010;
        25: y = 16'b0111111011101100;
        26: y = 16'b0111111110101010;
        27: y = 16'b0111111111111100;
        28: y = 16'b0111111111100000;
        29: y = 16'b0111111101011000;
        30: y = 16'b0111111001100100;
        31: y = 16'b0111110100000100;
        32: y = 16'b0111101100111010;
        33: y = 16'b0111100100001000;
        34: y = 16'b0111011001101110;
        35: y = 16'b0111001101101111;
        36: y = 16'b0111000000001111;
        37: y = 16'b0110110001001111;
        38: y = 16'b0110100000110011;
        39: y = 16'b0110001110111110;
        40: y = 16'b0101111011110100;
        41: y = 16'b0101100111011010;
        42: y = 16'b0101010001110100;
        43: y = 16'b0100111011000101;
        44: y = 16'b0100100011010100;
        45: y = 16'b0100001010100100;
        46: y = 16'b0011110000111100;
        47: y = 16'b0011010110100001;
        48: y = 16'b0010111011011000;
        49: y = 16'b0010011111100111;
        50: y = 16'b0010000011010101;
        51: y = 16'b0001100110100110;
        52: y = 16'b0001001001100010;
        53: y = 16'b0000101100001110;
        54: y = 16'b0000001110110000;
        55: y = 16'b1111110001010000;
        56: y = 16'b1111010011110010;
        57: y = 16'b1110110110011110;
        58: y = 16'b1110011001011010;
        59: y = 16'b1101111100101011;
        60: y = 16'b1101100000011001;
        61: y = 16'b1101000100101000;
        62: y = 16'b1100101001011111;
        63: y = 16'b1100001111000100;
        64: y = 16'b1011110101011100;
        65: y = 16'b1011011100101100;
        66: y = 16'b1011000100111011;
        67: y = 16'b1010101110001100;
        68: y = 16'b1010011000100110;
        69: y = 16'b1010000100001100;
        70: y = 16'b1001110001000010;
        71: y = 16'b1001011111001101;
        72: y = 16'b1001001110110001;
        73: y = 16'b1000111111110001;
        74: y = 16'b1000110010010001;
        75: y = 16'b1000100110010010;
        76: y = 16'b1000011011111000;
        77: y = 16'b1000010011000110;
        78: y = 16'b1000001011111100;
        79: y = 16'b1000000110011100;
        80: y = 16'b1000000010101000;
        81: y = 16'b1000000000100000;
        82: y = 16'b1000000000000100;
        83: y = 16'b1000000001010110;
        84: y = 16'b1000000100010100;
        85: y = 16'b1000001000111110;
        86: y = 16'b1000001111010011;
        87: y = 16'b1000010111010010;
        88: y = 16'b1000100000111001;
        89: y = 16'b1000101100000101;
        90: y = 16'b1000111000110101;
        91: y = 16'b1001000111000110;
        92: y = 16'b1001010110110100;
        93: y = 16'b1001100111111101;
        94: y = 16'b1001111010011100;
        95: y = 16'b1010001110001111;
        96: y = 16'b1010100011010000;
        97: y = 16'b1010111001011011;
        98: y = 16'b1011010000101100;
        99: y = 16'b1011101000111101;
        100: y = 16'b1100000010001001;
        101: y = 16'b1100011100001011;
        102: y = 16'b1100110110111110;
        103: y = 16'b1101010010011100;
        104: y = 16'b1101101110011110;
        105: y = 16'b1110001010111111;
        106: y = 16'b1110100111111010;
        107: y = 16'b1111000101000111;
        108: y = 16'b1111100010100000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=466.16Hz, Fs=48000Hz, 16-bit

module lut_As
(
    input      [6:0] x,
    output     [6:0] x_max,
    output reg [15:0] y
);

    assign x_max = 101;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011111100001;
        2: y = 16'b0000111110111011;
        3: y = 16'b0001011110000101;
        4: y = 16'b0001111100111000;
        5: y = 16'b0010011011001101;
        6: y = 16'b0010111000111101;
        7: y = 16'b0011010101111111;
        8: y = 16'b0011110010001110;
        9: y = 16'b0100001101100010;
        10: y = 16'b0100100111110100;
        11: y = 16'b0101000000111110;
        12: y = 16'b0101011000111011;
        13: y = 16'b0101101111100100;
        14: y = 16'b0110000100110011;
        15: y = 16'b0110011000100101;
        16: y = 16'b0110101010110011;
        17: y = 16'b0110111011011001;
        18: y = 16'b0111001010010100;
        19: y = 16'b0111010111011111;
        20: y = 16'b0111100010111000;
        21: y = 16'b0111101100011100;
        22: y = 16'b0111110100001000;
        23: y = 16'b0111111001111011;
        24: y = 16'b0111111101110011;
        25: y = 16'b0111111111101111;
        26: y = 16'b0111111111101111;
        27: y = 16'b0111111101110011;
        28: y = 16'b0111111001111011;
        29: y = 16'b0111110100001000;
        30: y = 16'b0111101100011100;
        31: y = 16'b0111100010111000;
        32: y = 16'b0111010111011111;
        33: y = 16'b0111001010010100;
        34: y = 16'b0110111011011001;
        35: y = 16'b0110101010110011;
        36: y = 16'b0110011000100101;
        37: y = 16'b0110000100110011;
        38: y = 16'b0101101111100100;
        39: y = 16'b0101011000111011;
        40: y = 16'b0101000000111110;
        41: y = 16'b0100100111110100;
        42: y = 16'b0100001101100010;
        43: y = 16'b0011110010001110;
        44: y = 16'b0011010101111111;
        45: y = 16'b0010111000111101;
        46: y = 16'b0010011011001101;
        47: y = 16'b0001111100111000;
        48: y = 16'b0001011110000101;
        49: y = 16'b0000111110111011;
        50: y = 16'b0000011111100001;
        51: y = 16'b0000000000000000;
        52: y = 16'b1111100000011111;
        53: y = 16'b1111000001000101;
        54: y = 16'b1110100001111011;
        55: y = 16'b1110000011001000;
        56: y = 16'b1101100100110011;
        57: y = 16'b1101000111000011;
        58: y = 16'b1100101010000001;
        59: y = 16'b1100001101110010;
        60: y = 16'b1011110010011110;
        61: y = 16'b1011011000001100;
        62: y = 16'b1010111111000010;
        63: y = 16'b1010100111000101;
        64: y = 16'b1010010000011100;
        65: y = 16'b1001111011001101;
        66: y = 16'b1001100111011011;
        67: y = 16'b1001010101001101;
        68: y = 16'b1001000100100111;
        69: y = 16'b1000110101101100;
        70: y = 16'b1000101000100001;
        71: y = 16'b1000011101001000;
        72: y = 16'b1000010011100100;
        73: y = 16'b1000001011111000;
        74: y = 16'b1000000110000101;
        75: y = 16'b1000000010001101;
        76: y = 16'b1000000000010001;
        77: y = 16'b1000000000010001;
        78: y = 16'b1000000010001101;
        79: y = 16'b1000000110000101;
        80: y = 16'b1000001011111000;
        81: y = 16'b1000010011100100;
        82: y = 16'b1000011101001000;
        83: y = 16'b1000101000100001;
        84: y = 16'b1000110101101100;
        85: y = 16'b1001000100100111;
        86: y = 16'b1001010101001101;
        87: y = 16'b1001100111011011;
        88: y = 16'b1001111011001101;
        89: y = 16'b1010010000011100;
        90: y = 16'b1010100111000101;
        91: y = 16'b1010111111000010;
        92: y = 16'b1011011000001100;
        93: y = 16'b1011110010011110;
        94: y = 16'b1100001101110010;
        95: y = 16'b1100101010000001;
        96: y = 16'b1101000111000011;
        97: y = 16'b1101100100110011;
        98: y = 16'b1110000011001000;
        99: y = 16'b1110100001111011;
        100: y = 16'b1111000001000101;
        101: y = 16'b1111100000011111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=493.88Hz, Fs=48000Hz, 16-bit

module lut_B
(
    input      [6:0] x,
    output     [6:0] x_max,
    output reg [15:0] y
);

    assign x_max = 96;

    always @ (*)
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000100001001001;
        2: y = 16'b0001000010001001;
        3: y = 16'b0001100010110111;
        4: y = 16'b0010000011001011;
        5: y = 16'b0010100010111100;
        6: y = 16'b0011000010000001;
        7: y = 16'b0011100000010010;
        8: y = 16'b0011111101100110;
        9: y = 16'b0100011001110111;
        10: y = 16'b0100110100111011;
        11: y = 16'b0101001110101101;
        12: y = 16'b0101100111000101;
        13: y = 16'b0101111101111101;
        14: y = 16'b0110010011001110;
        15: y = 16'b0110100110110011;
        16: y = 16'b0110111000100111;
        17: y = 16'b0111001000100100;
        18: y = 16'b0111010110100110;
        19: y = 16'b0111100010101010;
        20: y = 16'b0111101100101101;
        21: y = 16'b0111110100101100;
        22: y = 16'b0111111010100100;
        23: y = 16'b0111111110010100;
        24: y = 16'b0111111111111011;
        25: y = 16'b0111111111011000;
        26: y = 16'b0111111100101101;
        27: y = 16'b0111110111111001;
        28: y = 16'b0111110000111101;
        29: y = 16'b0111100111111100;
        30: y = 16'b0111011100111000;
        31: y = 16'b0111001111110101;
        32: y = 16'b0111000000110100;
        33: y = 16'b0110101111111011;
        34: y = 16'b0110011101001111;
        35: y = 16'b0110001000110011;
        36: y = 16'b0101110010101110;
        37: y = 16'b0101011011000101;
        38: y = 16'b0101000001111111;
        39: y = 16'b0100100111100011;
        40: y = 16'b0100001011110111;
        41: y = 16'b0011101111000100;
        42: y = 16'b0011010001010000;
        43: y = 16'b0010110010100100;
        44: y = 16'b0010010011001001;
        45: y = 16'b0001110011000101;
        46: y = 16'b0001010010100011;
        47: y = 16'b0000110001101011;
        48: y = 16'b0000010000100101;
        49: y = 16'b1111101111011011;
        50: y = 16'b1111001110010101;
        51: y = 16'b1110101101011101;
        52: y = 16'b1110001100111011;
        53: y = 16'b1101101100110111;
        54: y = 16'b1101001101011100;
        55: y = 16'b1100101110110000;
        56: y = 16'b1100010000111100;
        57: y = 16'b1011110100001001;
        58: y = 16'b1011011000011101;
        59: y = 16'b1010111110000001;
        60: y = 16'b1010100100111011;
        61: y = 16'b1010001101010010;
        62: y = 16'b1001110111001101;
        63: y = 16'b1001100010110001;
        64: y = 16'b1001010000000101;
        65: y = 16'b1000111111001100;
        66: y = 16'b1000110000001011;
        67: y = 16'b1000100011001000;
        68: y = 16'b1000011000000100;
        69: y = 16'b1000001111000011;
        70: y = 16'b1000001000000111;
        71: y = 16'b1000000011010011;
        72: y = 16'b1000000000101000;
        73: y = 16'b1000000000000101;
        74: y = 16'b1000000001101100;
        75: y = 16'b1000000101011100;
        76: y = 16'b1000001011010100;
        77: y = 16'b1000010011010011;
        78: y = 16'b1000011101010110;
        79: y = 16'b1000101001011010;
        80: y = 16'b1000110111011100;
        81: y = 16'b1001000111011001;
        82: y = 16'b1001011001001101;
        83: y = 16'b1001101100110010;
        84: y = 16'b1010000010000011;
        85: y = 16'b1010011000111011;
        86: y = 16'b1010110001010011;
        87: y = 16'b1011001011000101;
        88: y = 16'b1011100110001001;
        89: y = 16'b1100000010011010;
        90: y = 16'b1100011111101110;
        91: y = 16'b1100111101111111;
        92: y = 16'b1101011101000100;
        93: y = 16'b1101111100110101;
        94: y = 16'b1110011101001001;
        95: y = 16'b1110111101110111;
        96: y = 16'b1111011110110111;
        default: y = 16'b0;
        endcase

endmodule

