
`include "user_axis.sv"
`include "bind_user_axis.sv"
