// y(t) = sin(2*pi*F*t), F=1000Hz, Fs=48000Hz
0: y = 32'b00000000000000000000000000000000;
1: y = 32'b00010000101101010001010100001111;
2: y = 32'b00100001001000001111101110000011;
3: y = 32'b00110000111110111100010101001101;
4: y = 32'b00111111111111111111111111111111;
5: y = 32'b01001101111010111110010011111110;
6: y = 32'b01011010100000100111100110011001;
7: y = 32'b01100101100011001001101000101101;
8: y = 32'b01101110110110011110101110100001;
9: y = 32'b01110110010000011010111100111100;
10: y = 32'b01111011101000110111010100011100;
11: y = 32'b01111110111001111010101001001011;
12: y = 32'b01111111111111111111111111111111;
13: y = 32'b01111110111001111010101001001011;
14: y = 32'b01111011101000110111010100011100;
15: y = 32'b01110110010000011010111100111100;
16: y = 32'b01101110110110011110101110100001;
17: y = 32'b01100101100011001001101000101101;
18: y = 32'b01011010100000100111100110011001;
19: y = 32'b01001101111010111110010011111110;
20: y = 32'b00111111111111111111111111111111;
21: y = 32'b00110000111110111100010101001101;
22: y = 32'b00100001001000001111101110000011;
23: y = 32'b00010000101101010001010100001111;
24: y = 32'b00000000000000000000000000000000;
25: y = 32'b11101111010010101110101011110001;
26: y = 32'b11011110110111110000010001111101;
27: y = 32'b11001111000001000011101010110011;
28: y = 32'b11000000000000000000000000000001;
29: y = 32'b10110010000101000001101100000010;
30: y = 32'b10100101011111011000011001100111;
31: y = 32'b10011010011100110110010111010011;
32: y = 32'b10010001001001100001010001011111;
33: y = 32'b10001001101111100101000011000100;
34: y = 32'b10000100010111001000101011100100;
35: y = 32'b10000001000110000101010110110101;
36: y = 32'b10000000000000000000000000000001;
37: y = 32'b10000001000110000101010110110101;
38: y = 32'b10000100010111001000101011100100;
39: y = 32'b10001001101111100101000011000100;
40: y = 32'b10010001001001100001010001011111;
41: y = 32'b10011010011100110110010111010011;
42: y = 32'b10100101011111011000011001100111;
43: y = 32'b10110010000101000001101100000010;
44: y = 32'b11000000000000000000000000000000;
45: y = 32'b11001111000001000011101010110011;
46: y = 32'b11011110110111110000010001111101;
47: y = 32'b11101111010010101110101011110001;
