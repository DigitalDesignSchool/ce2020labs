
`include "bind_fifo_w8.sv"
`include "fifo_w8.sv"

