// This code on EDA Playground: https://edaplayground.com/x/kXW_

package riscv_instruction;

  // TODO parameters

  //--------------------------------------------------------------------------

  // TODO typedefs

  // TODO enums

  //--------------------------------------------------------------------------

  class riscv_instruction;

    // TODO rand fields

    //------------------------------------------------------------------------

    // TODO constraints

    //------------------------------------------------------------------------

    function string str ();

      string s;

      $sformat (s, "TODO fields");

      return s;

    endfunction

  endclass

endpackage
