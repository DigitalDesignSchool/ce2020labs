
`include "double_buffer.sv"
