
`include "skid_crd.sv"
 

