// Code your design here
module user();
  
  
endmodule