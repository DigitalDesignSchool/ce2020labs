
`include "fifo_256.sv"
`include "bind_fifo_256.sv"
