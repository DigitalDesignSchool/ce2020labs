`ifndef CONFIG_VH
`define CONFIG_VH

`timescale 1 ns / 1 ps

`endif
