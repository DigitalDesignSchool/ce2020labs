
`include "conv_with_fifo.sv"
`include "fifo_w8.sv" 
`include "ram256x16.sv"
