
`include "ram256x16.sv"
`include "ram256x256.sv"
`include "fifo_256.sv"
`include "credit_return.sv"
`include "binding_coverage_credit_return.sv"
