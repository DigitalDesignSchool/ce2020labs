`ifndef AXI_DEFINES
`define AXI_DEFINES

`define C_S00_BASEADDR 0
`define NO_OF_TRANSACTIONS 100
typedef enum {WRITE = 1, READ = 0} write_read_e;
`endif
