
`include "skid_buffer.sv"
 

